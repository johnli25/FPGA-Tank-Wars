module obstacle_array();





endmodule 